module TB (tb_CLK, tb_ENB, tb_DIR, tb_S_OUT, tb_)
